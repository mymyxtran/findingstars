`timescale 1ns/1ns

module draw_box();

endmodule

module drawDataPath(xLeft, xRight, yTop, yBottom, countXEn, countYEn, ld_x, ld_y, xEdge, yEdge, xOut, yOut, colOut);

	//these define the dimensions of the box
	input xLeft, xRight;
	input yTop, yBottom;
	
	

endmodule

module drawControl();

endmodule

