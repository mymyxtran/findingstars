`timescale 1ns/1ns

module clean_star();

endmodule

module cleanDataPath();



endmodule

module cleanControl();

endmodule

